module negador_1_bit (input logic a, output logic result);
										
	assign result = ~a;

endmodule 